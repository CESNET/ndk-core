//-- pkg.sv
//-- Copyright (C) 2023 CESNET z. s. p. o.
//-- Author(s): Daniel Kriz <danielkriz@cesnet.cz>

//-- SPDX-License-Identifier: BSD-3-Clause


`ifndef DOWN_HDR_PKG
`define DOWN_HDR_PKG

package uvm_down_hdr;

    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "tag_manager.sv"
    `include "sync_tag.sv"
    `include "config.sv"
    `include "sequence_item.sv"
    `include "sequence_item_dma_up.sv"
    `include "sequence_item_rq.sv"
    `include "sequencer.sv"
    `include "sequence.sv"
    `include "monitor.sv"
    `include "agent.sv"
    `include "encode_type.sv"

endpackage

`endif
